LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY FA IS PORT(
	A, B, D : in std_logic;
	S: out std_logic;
	C: out std_logic
);
END FA;

ARCHITECTURE BEHAVIORAL OF FA IS
BEGIN 

	C<= (A AND B)OR(B AND D)OR(A AND D);
	S<= A XOR B XOR D;

END BEHAVIORAL;