LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY HA IS PORT(
	A, B : in std_logic;
	S: out std_logic;
	C: out std_logic
);
END HA;

ARCHITECTURE BEHAVIORAL OF HA IS
BEGIN
	C<= A AND B;
	S<= A XOR B;

END BEHAVIORAL;
